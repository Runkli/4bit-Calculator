library verilog;
use verilog.vl_types.all;
entity ARS_vlg_vec_tst is
end ARS_vlg_vec_tst;
