library verilog;
use verilog.vl_types.all;
entity LRS_vlg_check_tst is
    port(
        Output          : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end LRS_vlg_check_tst;
