library verilog;
use verilog.vl_types.all;
entity LRS_vlg_vec_tst is
end LRS_vlg_vec_tst;
