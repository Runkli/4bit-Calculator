library verilog;
use verilog.vl_types.all;
entity LLS_vlg_vec_tst is
end LLS_vlg_vec_tst;
