library verilog;
use verilog.vl_types.all;
entity Calculator_vlg_vec_tst is
end Calculator_vlg_vec_tst;
