library verilog;
use verilog.vl_types.all;
entity LLS_vlg_check_tst is
    port(
        lls_out         : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end LLS_vlg_check_tst;
